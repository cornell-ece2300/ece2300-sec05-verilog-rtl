//========================================================================
// AbsDiff_4b_RTL
//========================================================================

`ifndef ABS_DIFF_4B_RTL_V
`define ABS_DIFF_4B_RTL_V

//''' ACTIVITY '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''
// Include any other hardware modules as necessary
//''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

module AbsDiff_4b_RTL
(
  (* keep=1 *) input  logic [3:0] in0,
  (* keep=1 *) input  logic [3:0] in1,
  (* keep=1 *) output logic [3:0] diff
);

  //''' ACTIVITY '''''''''''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement 4b absolute difference unit using RTL
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

`endif /* ABS_DIFF_4B_RTL_V */
