//========================================================================
// Mux2_4b_RTL
//========================================================================

`ifndef MUX2_4B_RTL
`define MUX2_4B_RTL

module Mux2_4b_RTL
(
  (* keep=1 *) input  logic [3:0] in0,
  (* keep=1 *) input  logic [3:0] in1,
  (* keep=1 *) input  logic       sel,
  (* keep=1 *) output logic [3:0] out
);

  //''' ACTIVITY '''''''''''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement 4b mux using RTL
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

`endif /* MUX2_4B_RTL */

